
	parameter WB_ADDR_WIDTH = 2;	
	parameter WB_DATA_WIDTH = 8;

